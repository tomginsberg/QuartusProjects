-- jtag_io.vhd

-- Generated using ACDS version 15.0 150

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity jtag_io is
	port (
		tms : in  std_logic := '0'; -- jtag.tms
		tdi : in  std_logic := '0'; --     .tdi
		tdo : out std_logic;        --     .tdo
		tck : in  std_logic := '0'  --  tck.clk
	);
end entity jtag_io;

architecture rtl of jtag_io is
	component altera_soft_core_jtag_io is
		generic (
			ENABLE_JTAG_IO_SELECTION : integer := 0
		);
		port (
			tms         : in  std_logic := 'X'; -- tms
			tdi         : in  std_logic := 'X'; -- tdi
			tdo         : out std_logic;        -- tdo
			tck         : in  std_logic := 'X'; -- clk
			select_this : in  std_logic := 'X'  -- select_this
		);
	end component altera_soft_core_jtag_io;

begin

	jtag_io_inst : component altera_soft_core_jtag_io
		generic map (
			ENABLE_JTAG_IO_SELECTION => 0
		)
		port map (
			tms         => tms, -- jtag.tms
			tdi         => tdi, --     .tdi
			tdo         => tdo, --     .tdo
			tck         => tck, --  tck.clk
			select_this => '0'  -- (terminated)
		);

end architecture rtl; -- of jtag_io
